package spi_pkg;
//`include "interface.sv"
import uvm_pkg::*;
`include "uvm_macros.svh"
`include "spi_sequence_item.sv"
`include "spi_sequence.sv"
`include "spi_sequence2.sv"
`include "spi_sequence3.sv"
`include "spi_sequence4.sv"
`include "spi_sequence5.sv"
`include "spi_sequence6.sv"
`include "spi_driver.sv"
`include "spi_sequencer.sv"
`include "spi_virtual_sequencer.sv"
`include "spi_virtual_sequence.sv"
`include "spi_scoreboard.sv"
`include "collector.sv"
`include "spi_monitor.sv"
`include "spi_agent.sv"
`include "spi_environment.sv"
`include "spi_test.sv"

endpackage